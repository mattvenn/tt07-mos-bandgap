magic
tech sky130A
magscale 1 2
timestamp 1716715833
<< nwell >>
rect 1420 740 1480 1040
<< viali >>
rect 40 3600 200 3660
rect 740 3600 900 3660
rect 1440 3600 1600 3660
rect 20 2020 200 2080
rect 720 2020 900 2080
rect 20 1100 200 1160
rect 720 1100 900 1160
rect 1420 1100 1600 1160
rect -680 620 -460 680
rect 2120 620 2340 680
<< metal1 >>
rect -800 3900 2400 4200
rect -600 3440 -520 3446
rect -600 3354 -520 3360
rect -300 1300 -160 3900
rect -100 3860 1720 3900
rect -100 3780 1060 3860
rect 1140 3780 1720 3860
rect -100 3660 1720 3780
rect -100 3600 40 3660
rect 200 3600 740 3660
rect 900 3600 1440 3660
rect 1600 3600 1720 3660
rect -100 3440 0 3600
rect 28 3594 212 3600
rect 728 3594 912 3600
rect 1428 3594 1612 3600
rect 80 3480 1560 3560
rect -100 3240 80 3440
rect 140 3060 200 3440
rect 400 3060 480 3480
rect 1640 3440 1720 3600
rect 2180 3440 2760 3540
rect 140 2980 480 3060
rect 0 2860 80 2866
rect 0 2220 80 2780
rect 140 2220 200 2980
rect 720 2760 780 3440
rect 1040 3400 1160 3420
rect 840 3320 1060 3400
rect 1140 3320 1160 3400
rect 1040 3300 1160 3320
rect 1420 2980 1480 3440
rect 1540 3240 1720 3440
rect 1820 3360 2760 3440
rect 1820 2980 1900 3360
rect 2180 3280 2760 3360
rect 1420 2900 1900 2980
rect 420 2700 780 2760
rect 420 2180 480 2700
rect 720 2220 780 2700
rect 840 2220 1120 2420
rect 80 2120 860 2180
rect 8 2080 212 2086
rect 708 2080 912 2086
rect -80 2020 20 2080
rect 200 2020 720 2080
rect 900 2020 980 2080
rect -80 2000 980 2020
rect 360 1840 560 2000
rect 340 1820 580 1840
rect 340 1620 360 1820
rect 560 1620 580 1820
rect 340 1600 580 1620
rect 1060 1430 1120 2220
rect 1060 1360 1120 1370
rect -300 1160 1720 1300
rect -300 1100 20 1160
rect 200 1100 720 1160
rect 900 1100 1420 1160
rect 1600 1100 1720 1160
rect 8 1094 212 1100
rect 708 1094 912 1100
rect 1408 1094 1612 1100
rect -620 840 80 1020
rect 140 840 360 1020
rect 354 820 360 840
rect 560 840 780 1020
rect 840 950 1120 1020
rect 840 890 1060 950
rect 1120 890 1126 950
rect 840 840 1120 890
rect 560 820 566 840
rect 360 780 560 820
rect 1420 780 1480 1040
rect 1540 840 2280 1020
rect 80 700 860 780
rect -780 680 -340 700
rect -780 620 -680 680
rect -460 620 -340 680
rect -780 500 -340 620
rect 360 500 560 700
rect 1420 500 1600 780
rect 2108 680 2352 686
rect 2000 620 2120 680
rect 2340 620 2400 680
rect 2000 500 2400 620
rect -800 200 2400 500
<< via1 >>
rect -600 3360 -520 3440
rect 1060 3780 1140 3860
rect 0 2780 80 2860
rect 1060 3320 1140 3400
rect 360 1620 560 1820
rect 1060 1370 1120 1430
rect 360 820 560 1020
rect 1060 890 1120 950
<< metal2 >>
rect 1040 3860 1160 3880
rect 1040 3780 1060 3860
rect 1140 3780 1160 3860
rect -606 3360 -600 3440
rect -520 3360 -360 3440
rect -440 2860 -360 3360
rect 1040 3400 1160 3780
rect 1040 3320 1060 3400
rect 1140 3320 1160 3400
rect 1040 3300 1160 3320
rect -440 2780 0 2860
rect 80 2780 86 2860
rect 340 1820 580 1840
rect 340 1620 360 1820
rect 560 1620 580 1820
rect 340 1600 580 1620
rect 360 1020 560 1600
rect 1054 1370 1060 1430
rect 1120 1370 1126 1430
rect 1060 950 1120 1370
rect 1060 884 1120 890
rect 360 814 560 820
use sky130_fd_pr__pfet_01v8_MGS3BN  XM1
timestamp 1716712743
transform 1 0 111 0 1 3384
box -211 -284 211 284
use sky130_fd_pr__pfet_01v8_MGS3BN  XM2
timestamp 1716712743
transform 1 0 811 0 1 3384
box -211 -284 211 284
use sky130_fd_pr__pfet_01v8_MGS3BN  XM3
timestamp 1716712743
transform 1 0 1511 0 1 3384
box -211 -284 211 284
use sky130_fd_pr__nfet_01v8_64QSBY  XM4
timestamp 1716713073
transform 1 0 111 0 1 2279
box -211 -279 211 279
use sky130_fd_pr__nfet_01v8_64QSBY  XM5
timestamp 1716713073
transform 1 0 811 0 1 2279
box -211 -279 211 279
use sky130_fd_pr__pfet_01v8_LGS3BL  XM6
timestamp 1716713827
transform 1 0 111 0 1 884
box -211 -284 211 284
use sky130_fd_pr__pfet_01v8_LGS3BL  XM7
timestamp 1716713827
transform 1 0 811 0 1 884
box -211 -284 211 284
use sky130_fd_pr__pfet_01v8_LGS3BL  XM8
timestamp 1716713827
transform 1 0 1511 0 1 884
box -211 -284 211 284
use sky130_fd_pr__res_high_po_0p69_CY6CB8  XR1
timestamp 1716712743
transform 1 0 2235 0 1 2182
box -235 -1582 235 1582
use sky130_fd_pr__res_high_po_0p69_CY6CB8  XR4
timestamp 1716712743
transform 1 0 -565 0 1 2182
box -235 -1582 235 1582
<< labels >>
flabel metal1 2100 4000 2300 4200 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal1 2100 300 2300 500 0 FreeSans 256 0 0 0 VSS
port 2 nsew
flabel metal1 2560 3320 2760 3520 0 FreeSans 256 0 0 0 vref
port 1 nsew
flabel metal2 -440 2780 0 2860 0 FreeSans 800 0 0 0 Va
flabel space 1060 840 1120 2420 0 FreeSans 800 0 0 0 Vb
flabel metal1 140 2980 480 3060 0 FreeSans 800 0 0 0 top_gate
flabel metal1 420 2700 780 2760 0 FreeSans 800 0 0 0 n_gate
flabel metal1 1540 840 2280 1020 0 FreeSans 800 0 0 0 r1_m8
flabel metal1 -620 840 80 1020 0 FreeSans 800 0 0 0 r4_m6
<< end >>
