magic
tech sky130A
magscale 1 2
timestamp 1716717956
<< metal1 >>
rect 18050 12990 18350 12996
rect 18350 12690 26050 12990
rect 18050 12684 18350 12690
rect 21150 7050 21450 12690
rect 30530 12210 30750 12216
rect 28450 11990 30530 12210
rect 30530 11984 30750 11990
rect 23110 9210 23410 9216
rect 23410 8910 25930 9210
rect 23110 8904 23410 8910
rect 21150 6750 25890 7050
rect 23590 2410 23890 2416
rect 23890 2110 25850 2410
rect 23590 2104 23890 2110
<< via1 >>
rect 18050 12690 18350 12990
rect 30530 11990 30750 12210
rect 23110 8910 23410 9210
rect 23590 2110 23890 2410
<< metal2 >>
rect 11875 12990 12165 12994
rect 11870 12985 18050 12990
rect 11870 12695 11875 12985
rect 12165 12695 18050 12985
rect 11870 12690 18050 12695
rect 18350 12690 18356 12990
rect 11875 12686 12165 12690
rect 30524 11990 30530 12210
rect 30750 11990 30756 12210
rect 22015 9210 22305 9214
rect 22010 9205 23110 9210
rect 22010 8915 22015 9205
rect 22305 8915 23110 9205
rect 22010 8910 23110 8915
rect 23410 8910 23416 9210
rect 22015 8906 22305 8910
rect 29560 6420 29960 6430
rect 29560 6050 29960 6060
rect 30530 5345 30750 11990
rect 30526 5135 30535 5345
rect 30745 5135 30754 5345
rect 30530 5130 30750 5135
rect 26380 3440 26540 3450
rect 28400 3420 28540 3430
rect 28400 3290 28540 3300
rect 26380 3270 26540 3280
rect 21855 2410 22145 2414
rect 21850 2405 23590 2410
rect 21850 2115 21855 2405
rect 22145 2115 23590 2405
rect 21850 2110 23590 2115
rect 23890 2110 23896 2410
rect 21855 2106 22145 2110
<< via2 >>
rect 11875 12695 12165 12985
rect 22015 8915 22305 9205
rect 29560 6060 29960 6420
rect 30535 5135 30745 5345
rect 26380 3280 26540 3440
rect 28400 3300 28540 3420
rect 21855 2115 22145 2405
<< metal3 >>
rect 6431 12990 6729 12995
rect 6430 12989 12170 12990
rect 6430 12691 6431 12989
rect 6729 12985 12170 12989
rect 6729 12695 11875 12985
rect 12165 12695 12170 12985
rect 6729 12691 12170 12695
rect 6430 12690 12170 12691
rect 6431 12685 6729 12690
rect 20551 9210 20849 9215
rect 20550 9209 22310 9210
rect 20550 8911 20551 9209
rect 20849 9205 22310 9209
rect 20849 8915 22015 9205
rect 22305 8915 22310 9205
rect 20849 8911 22310 8915
rect 20550 8910 22310 8911
rect 20551 8905 20849 8910
rect 29480 6420 30980 6440
rect 29480 6120 29560 6420
rect 29550 6060 29560 6120
rect 29960 6350 30980 6420
rect 31283 6350 31461 6355
rect 29960 6349 31462 6350
rect 29960 6171 31283 6349
rect 31461 6171 31462 6349
rect 29960 6170 31462 6171
rect 29960 6120 30980 6170
rect 31283 6165 31461 6170
rect 29960 6060 29970 6120
rect 29550 6055 29970 6060
rect 30530 5345 30750 5350
rect 30530 5135 30535 5345
rect 30745 5135 30750 5345
rect 24740 3440 26600 3520
rect 30530 3480 30750 5135
rect 24740 3280 26380 3440
rect 26540 3280 26600 3440
rect 28360 3420 30750 3480
rect 28360 3300 28400 3420
rect 28540 3300 30750 3420
rect 19991 2410 20289 2415
rect 19990 2409 22150 2410
rect 19990 2111 19991 2409
rect 20289 2405 22150 2409
rect 20289 2115 21855 2405
rect 22145 2115 22150 2405
rect 20289 2111 22150 2115
rect 19990 2110 22150 2111
rect 19991 2105 20289 2110
rect 24760 1740 25000 3280
rect 26370 3275 26550 3280
rect 28360 3260 30750 3300
rect 24760 1500 30500 1740
rect 30740 1500 30746 1740
<< via3 >>
rect 6431 12691 6729 12989
rect 20551 8911 20849 9209
rect 31283 6171 31461 6349
rect 19991 2111 20289 2409
rect 30500 1500 30740 1740
<< metal4 >>
rect 798 44770 858 45152
rect 1534 44770 1594 45152
rect 2270 44770 2330 45152
rect 3006 44770 3066 45152
rect 3742 44770 3802 45152
rect 4478 44770 4538 45152
rect 5214 44770 5274 45152
rect 5950 44770 6010 45152
rect 6686 44770 6746 45152
rect 7422 44770 7482 45152
rect 8158 44770 8218 45152
rect 8894 44770 8954 45152
rect 9630 44770 9690 45152
rect 10366 44770 10426 45152
rect 11102 44770 11162 45152
rect 11838 44770 11898 45152
rect 12574 44770 12634 45152
rect 13310 44770 13370 45152
rect 14046 44770 14106 45152
rect 14782 44770 14842 45152
rect 15518 44770 15578 45152
rect 16254 44770 16314 45152
rect 16990 44770 17050 45152
rect 17726 44770 17786 45152
rect 18462 44952 18522 45152
rect 19198 44952 19258 45152
rect 19934 44952 19994 45152
rect 20670 44952 20730 45152
rect 21406 44952 21466 45152
rect 22142 44952 22202 45152
rect 22878 44952 22938 45152
rect 23614 44952 23674 45152
rect 24350 44952 24410 45152
rect 25086 44952 25146 45152
rect 25822 44952 25882 45152
rect 26558 44952 26618 45152
rect 27294 44952 27354 45152
rect 28030 44952 28090 45152
rect 28766 44952 28826 45152
rect 29502 44952 29562 45152
rect 30238 44952 30298 45152
rect 30974 44952 31034 45152
rect 31710 44952 31770 45152
rect 570 44710 17786 44770
rect 9930 44152 9990 44710
rect 200 12990 500 44152
rect 200 12989 6730 12990
rect 200 12691 6431 12989
rect 6729 12691 6730 12989
rect 200 12690 6730 12691
rect 200 1000 500 12690
rect 9800 9210 10100 44152
rect 9800 9209 20850 9210
rect 9800 8911 20551 9209
rect 20849 8911 20850 9209
rect 9800 8910 20850 8911
rect 9800 1000 10100 8910
rect 19990 2409 20290 8910
rect 19990 2111 19991 2409
rect 20289 2111 20290 2409
rect 19990 2110 20290 2111
rect 31282 6349 31462 6350
rect 31282 6171 31283 6349
rect 31461 6171 31462 6349
rect 30499 1740 30741 1741
rect 31282 1740 31462 6171
rect 30499 1500 30500 1740
rect 30740 1500 31462 1740
rect 30499 1499 30741 1500
rect 370 0 550 200
rect 4786 0 4966 200
rect 9202 0 9382 200
rect 13618 0 13798 200
rect 18034 0 18214 200
rect 22450 0 22630 200
rect 26866 0 27046 200
rect 31282 0 31462 1500
use bandgap  bandgap_0
timestamp 1716715833
transform 1 0 25990 0 1 8722
box -800 200 2760 4200
use p3_opamp  p3_opamp_0
timestamp 1715778954
transform 1 0 21684 0 1 -1096
box 3650 3170 8500 8260
<< labels >>
flabel metal4 s 30974 44952 31034 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 31710 44952 31770 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 30238 44952 30298 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 31282 0 31462 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26866 0 27046 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22450 0 22630 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18034 0 18214 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 13618 0 13798 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 9202 0 9382 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 4786 0 4966 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 370 0 550 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 29502 44952 29562 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 28030 44952 28090 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 27294 44952 27354 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 25822 44952 25882 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 25086 44952 25146 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23614 44952 23674 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22878 44952 22938 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21406 44952 21466 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 20670 44952 20730 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19198 44952 19258 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 18462 44952 18522 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 5950 44952 6010 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 5214 44952 5274 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 4478 44952 4538 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 3742 44952 3802 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 3006 44952 3066 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 2270 44952 2330 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 1534 44952 1594 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 798 44952 858 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 11838 44952 11898 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 10366 44952 10426 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 9630 44952 9690 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 8158 44952 8218 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 7422 44952 7482 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 16990 44952 17050 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 16254 44952 16314 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 14782 44952 14842 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 14046 44952 14106 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 12574 44952 12634 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 500 44152 1 FreeSans 4800 0 0 0 VPWR
port 51 nsew power bidirectional
flabel metal4 9800 1000 10100 44152 1 FreeSans 4800 0 0 0 VGND
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
