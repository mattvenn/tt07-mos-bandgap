magic
tech sky130A
magscale 1 2
timestamp 1717066714
<< viali >>
rect 1000 8400 1080 10260
rect 3800 8420 3900 10200
rect 6620 8420 6700 10260
rect -1842 5756 -1686 6210
rect 280 5780 400 6180
rect 9580 5780 9680 6180
rect 11680 5780 11800 6180
rect -1080 5620 -480 5680
rect 10420 5600 10960 5700
rect 2000 5420 3020 5480
rect 4800 5400 5740 5480
rect 2160 4880 2940 5000
rect 6880 4880 7480 4940
rect 4800 3620 5320 3700
<< metal1 >>
rect -2000 11940 11800 12200
rect -2000 11440 8240 11940
rect 8740 11440 11800 11940
rect -2000 11200 11800 11440
rect 860 10300 1000 11200
rect 1220 10680 3520 10700
rect 1220 10440 2020 10680
rect 2360 10440 3520 10680
rect 1220 10380 3520 10440
rect 860 10260 1200 10300
rect 860 8400 1000 10260
rect 1080 8400 1200 10260
rect 860 8380 1200 8400
rect 3200 8360 3520 10380
rect 3660 10300 3800 11200
rect 4020 10680 6000 10700
rect 4020 10440 4820 10680
rect 5160 10440 6000 10680
rect 4020 10380 6000 10440
rect 3660 10200 4000 10300
rect 3660 8420 3800 10200
rect 3900 8420 4000 10200
rect 3660 8380 4000 8420
rect 6000 8360 6280 10340
rect 6460 10300 6600 11200
rect 6820 10680 8800 10700
rect 6820 10440 7640 10680
rect 7980 10440 8800 10680
rect 6820 10380 8800 10440
rect 6460 10260 6800 10300
rect 6460 8420 6620 10260
rect 6700 8420 6800 10260
rect 6460 8380 6800 8420
rect 8800 8360 9280 10320
rect 2020 7880 2980 7940
rect 2020 7660 2320 7880
rect 2660 7660 2980 7880
rect 2020 7580 2980 7660
rect 3380 7540 3520 8360
rect 6140 7940 6280 8360
rect 4620 7880 6280 7940
rect 4620 7660 4940 7880
rect 5280 7660 6280 7880
rect 4620 7620 6280 7660
rect 4620 7580 5860 7620
rect -1860 6210 -1660 6240
rect -1860 5756 -1842 6210
rect -1686 5756 -1660 6210
rect 1520 6200 1980 7540
rect 260 6180 1980 6200
rect 260 5780 280 6180
rect 400 5780 1980 6180
rect 260 5760 1980 5780
rect -1860 4740 -1660 5756
rect -1110 5600 -1100 5700
rect -460 5600 -450 5700
rect 1520 5560 1980 5760
rect 3000 7400 3520 7540
rect 3000 5560 3260 7400
rect 1980 5480 3080 5500
rect 1980 5420 2000 5480
rect 3020 5420 3080 5480
rect 1980 5360 3080 5420
rect 1980 5240 3280 5360
rect 2130 4860 2140 5020
rect 2960 4860 2970 5020
rect 3160 4820 3280 5240
rect -1860 4100 2000 4740
rect 1720 2880 2000 4100
rect 3000 2780 3280 4820
rect 4480 3700 4601 7360
rect 5600 5560 5860 7580
rect 9040 7460 9280 8360
rect 8000 6200 9280 7460
rect 8000 6180 9700 6200
rect 8000 5780 9580 6180
rect 9680 5780 9700 6180
rect 9040 5760 9700 5780
rect 11640 6180 11880 6220
rect 11640 5780 11680 6180
rect 11800 5780 11880 6180
rect 9040 5740 9280 5760
rect 10390 5560 10400 5740
rect 10980 5560 10990 5740
rect 4780 5480 5780 5500
rect 4780 5400 4800 5480
rect 5740 5400 5780 5480
rect 4780 5280 5780 5400
rect 4480 2960 4600 3700
rect 4770 3600 4780 3720
rect 5340 3600 5350 3720
rect 5660 3560 5780 5280
rect 6850 4840 6860 4980
rect 7480 4946 7490 4980
rect 7480 4874 7492 4946
rect 7480 4840 7490 4874
rect 5560 2920 5780 3560
rect 4720 2780 5780 2920
rect 6560 2780 6800 4820
rect 11640 4760 11880 5780
rect 7800 4380 11880 4760
rect 7800 2820 7980 4380
rect 2060 2760 6800 2780
rect 6880 2760 7720 2780
rect 2060 2560 7720 2760
rect 2000 2420 7720 2560
rect 2000 2000 7800 2420
rect -2000 1760 11800 2000
rect -2000 1320 -1100 1760
rect -460 1700 11800 1760
rect -460 1320 10420 1700
rect 10960 1320 11800 1700
rect -2000 1000 11800 1320
<< via1 >>
rect 8240 11440 8740 11940
rect 2020 10440 2360 10680
rect 4820 10440 5160 10680
rect 7640 10440 7980 10680
rect 2320 7660 2660 7880
rect 4940 7660 5280 7880
rect -1100 5680 -460 5700
rect -1100 5620 -1080 5680
rect -1080 5620 -480 5680
rect -480 5620 -460 5680
rect -1100 5600 -460 5620
rect 2140 5000 2960 5020
rect 2140 4880 2160 5000
rect 2160 4880 2940 5000
rect 2940 4880 2960 5000
rect 2140 4860 2960 4880
rect 10400 5700 10980 5740
rect 10400 5600 10420 5700
rect 10420 5600 10960 5700
rect 10960 5600 10980 5700
rect 10400 5560 10980 5600
rect 4780 3700 5340 3720
rect 4780 3620 4800 3700
rect 4800 3620 5320 3700
rect 5320 3620 5340 3700
rect 4780 3600 5340 3620
rect 6860 4940 7480 4980
rect 6860 4880 6880 4940
rect 6880 4880 7480 4940
rect 6860 4840 7480 4880
rect -1100 1320 -460 1760
rect 10420 1320 10960 1700
<< metal2 >>
rect 8180 11940 8780 12040
rect 8180 11440 8240 11940
rect 8740 11440 8780 11940
rect 2000 10680 8000 10720
rect 2000 10440 2020 10680
rect 2360 10440 4820 10680
rect 5160 10440 7640 10680
rect 7980 10440 8000 10680
rect 2000 10420 8000 10440
rect 8180 8920 8780 11440
rect 6900 8320 8780 8920
rect 2300 7880 5300 7900
rect 2300 7660 2320 7880
rect 2660 7660 4940 7880
rect 5280 7660 5300 7880
rect 2300 7640 5300 7660
rect -1140 5700 -420 5740
rect -1140 5600 -1100 5700
rect -460 5600 -420 5700
rect -1140 1760 -420 5600
rect 6900 5220 7500 8320
rect 2060 5020 7500 5220
rect 2060 4860 2140 5020
rect 2960 4980 7500 5020
rect 2960 4860 6860 4980
rect 2060 4840 6860 4860
rect 7480 4840 7500 4980
rect 2060 4620 7500 4840
rect 10380 5740 11000 5820
rect 10380 5560 10400 5740
rect 10980 5560 11000 5740
rect 4760 3720 5360 4620
rect 4760 3600 4780 3720
rect 5340 3600 5360 3720
rect 4760 3500 5360 3600
rect -1140 1320 -1100 1760
rect -460 1320 -420 1760
rect -1140 1260 -420 1320
rect 10380 1700 11000 5560
rect 10380 1320 10420 1700
rect 10960 1320 11000 1700
rect 10380 1280 11000 1320
use sky130_fd_pr__pfet_01v8_XLZ98A  XM1
timestamp 1717064607
transform 1 0 2196 0 1 9384
box -1196 -1184 1196 1184
use sky130_fd_pr__pfet_01v8_XLZ98A  XM2
timestamp 1717064607
transform 1 0 4996 0 1 9384
box -1196 -1184 1196 1184
use sky130_fd_pr__pfet_01v8_XLZ98A  XM3
timestamp 1717064607
transform 1 0 7796 0 1 9384
box -1196 -1184 1196 1184
use sky130_fd_pr__nfet_01v8_lvt_QYU87T  XM4
timestamp 1717064607
transform 1 0 5096 0 1 6579
box -696 -1179 696 1179
use sky130_fd_pr__pfet_01v8_lvt_GUWLND  XM5
timestamp 1717065751
transform 1 0 2496 0 1 3784
box -696 -1184 696 1184
use sky130_fd_pr__pfet_01v8_lvt_GUWLND  XM6
timestamp 1717065751
transform 1 0 7296 0 1 3784
box -696 -1184 696 1184
use sky130_fd_pr__pfet_01v8_lvt_3VXSVM  XM7
timestamp 1717065751
transform 1 0 5076 0 1 3224
box -696 -484 696 484
use sky130_fd_pr__nfet_01v8_lvt_QYU87T  XM9
timestamp 1717064607
transform 1 0 2496 0 1 6579
box -696 -1179 696 1179
use sky130_fd_pr__res_high_po_0p69_77P8PF  XR1
timestamp 1717064607
transform 1 0 10688 0 1 8084
box -1288 -2484 1288 2484
use sky130_fd_pr__res_high_po_0p69_77P8PF  XR4
timestamp 1717064607
transform 1 0 -712 0 1 8084
box -1288 -2484 1288 2484
<< labels >>
flabel metal1 -2000 11200 11800 12200 0 FreeSans 1600 0 0 0 VDD
port 3 nsew
flabel metal1 -2000 1000 11800 2000 0 FreeSans 1600 0 0 0 VSS
port 2 nsew
flabel metal2 2360 10420 4820 10720 0 FreeSans 1600 0 0 0 top_gate
flabel metal2 2660 7640 4940 7900 0 FreeSans 1600 0 0 0 n_gate
flabel metal1 8000 5780 9280 7460 0 FreeSans 1600 0 0 0 vref
port 4 nsew
flabel metal1 400 5760 1980 6200 0 FreeSans 1600 0 0 0 Va
flabel metal1 -1860 4100 1740 4740 0 FreeSans 1600 0 0 0 r4_m6
flabel metal1 7800 4380 11880 4760 0 FreeSans 1600 0 0 0 r1_m8
flabel metal1 4480 3700 4601 7360 0 FreeSans 1600 0 0 0 Vb
<< end >>
