magic
tech sky130A
magscale 1 2
timestamp 1717164048
<< metal1 >>
rect 15866 42828 16166 42834
rect 16166 42528 18040 42828
rect 15866 42522 16166 42528
rect 27846 36946 28066 37658
rect 27840 36726 27846 36946
rect 28066 36726 28072 36946
rect 22194 31008 22494 31014
rect 22582 31008 22882 32268
rect 22494 30708 22882 31008
rect 22194 30702 22494 30708
rect 20916 28868 21216 28874
rect 21216 28848 22540 28868
rect 21216 28568 25890 28848
rect 20916 28562 21216 28568
rect 22222 28548 25890 28568
rect 23590 24208 23890 24214
rect 23890 23908 25850 24208
rect 23590 23902 23890 23908
rect 15866 21030 16166 21036
rect 16166 20730 18040 21030
rect 15866 20724 16166 20730
rect 27846 15148 28066 15860
rect 27840 14928 27846 15148
rect 28066 14928 28072 15148
rect 22194 9210 22494 9216
rect 22582 9210 22882 10470
rect 22494 8910 22882 9210
rect 22194 8904 22494 8910
rect 20916 7070 21216 7076
rect 21216 7050 22540 7070
rect 21216 6770 25890 7050
rect 20916 6764 21216 6770
rect 22222 6750 25890 6770
rect 23590 2410 23890 2416
rect 23890 2110 25850 2410
rect 23590 2104 23890 2110
<< via1 >>
rect 15866 42528 16166 42828
rect 27846 36726 28066 36946
rect 22194 30708 22494 31008
rect 20916 28568 21216 28868
rect 23590 23908 23890 24208
rect 15866 20730 16166 21030
rect 27846 14928 28066 15148
rect 22194 8910 22494 9210
rect 20916 6770 21216 7070
rect 23590 2110 23890 2410
<< metal2 >>
rect 15001 42828 15291 42832
rect 14996 42823 15866 42828
rect 14996 42533 15001 42823
rect 15291 42533 15866 42823
rect 14996 42528 15866 42533
rect 16166 42528 16172 42828
rect 15001 42524 15291 42528
rect 27846 36946 28066 36952
rect 21583 31008 21873 31012
rect 21578 31003 22194 31008
rect 21578 30713 21583 31003
rect 21873 30713 22194 31003
rect 21578 30708 22194 30713
rect 22494 30708 22500 31008
rect 27846 30852 28066 36726
rect 21583 30704 21873 30708
rect 27846 30632 30750 30852
rect 20511 28868 20801 28872
rect 20506 28863 20916 28868
rect 20506 28573 20511 28863
rect 20801 28573 20916 28863
rect 20506 28568 20916 28573
rect 21216 28568 21222 28868
rect 20511 28564 20801 28568
rect 29560 28218 29960 28228
rect 29560 27848 29960 27858
rect 30530 27143 30750 30632
rect 30526 26933 30535 27143
rect 30745 26933 30754 27143
rect 30530 26928 30750 26933
rect 26380 25238 26540 25248
rect 28400 25218 28540 25228
rect 28400 25088 28540 25098
rect 26380 25068 26540 25078
rect 21855 24208 22145 24212
rect 21850 24203 23590 24208
rect 21850 23913 21855 24203
rect 22145 23913 23590 24203
rect 21850 23908 23590 23913
rect 23890 23908 23896 24208
rect 21855 23904 22145 23908
rect 15001 21030 15291 21034
rect 14996 21025 15866 21030
rect 14996 20735 15001 21025
rect 15291 20735 15866 21025
rect 14996 20730 15866 20735
rect 16166 20730 16172 21030
rect 15001 20726 15291 20730
rect 27846 15148 28066 15154
rect 21583 9210 21873 9214
rect 21578 9205 22194 9210
rect 21578 8915 21583 9205
rect 21873 8915 22194 9205
rect 21578 8910 22194 8915
rect 22494 8910 22500 9210
rect 27846 9054 28066 14928
rect 21583 8906 21873 8910
rect 27846 8834 30750 9054
rect 20511 7070 20801 7074
rect 20506 7065 20916 7070
rect 20506 6775 20511 7065
rect 20801 6775 20916 7065
rect 20506 6770 20916 6775
rect 21216 6770 21222 7070
rect 20511 6766 20801 6770
rect 29560 6420 29960 6430
rect 29560 6050 29960 6060
rect 30530 5345 30750 8834
rect 30526 5135 30535 5345
rect 30745 5135 30754 5345
rect 30530 5130 30750 5135
rect 26380 3440 26540 3450
rect 28400 3420 28540 3430
rect 28400 3290 28540 3300
rect 26380 3270 26540 3280
rect 21855 2410 22145 2414
rect 21850 2405 23590 2410
rect 21850 2115 21855 2405
rect 22145 2115 23590 2405
rect 21850 2110 23590 2115
rect 23890 2110 23896 2410
rect 21855 2106 22145 2110
<< via2 >>
rect 15001 42533 15291 42823
rect 21583 30713 21873 31003
rect 20511 28573 20801 28863
rect 29560 27858 29960 28218
rect 30535 26933 30745 27143
rect 26380 25078 26540 25238
rect 28400 25098 28540 25218
rect 21855 23913 22145 24203
rect 15001 20735 15291 21025
rect 21583 8915 21873 9205
rect 20511 6775 20801 7065
rect 29560 6060 29960 6420
rect 30535 5135 30745 5345
rect 26380 3280 26540 3440
rect 28400 3300 28540 3420
rect 21855 2115 22145 2405
<< metal3 >>
rect 12998 42823 15296 42828
rect 12998 42533 15001 42823
rect 15291 42533 15296 42823
rect 12998 42528 15296 42533
rect 12998 34788 13298 42528
rect 4766 34488 4772 34788
rect 5072 34488 13298 34788
rect 12998 28868 13298 34488
rect 20895 31008 21193 31013
rect 20894 31007 21878 31008
rect 20894 30709 20895 31007
rect 21193 31003 21878 31007
rect 21193 30713 21583 31003
rect 21873 30713 21878 31003
rect 21193 30709 21878 30713
rect 20894 30708 21878 30709
rect 20895 30703 21193 30708
rect 12998 28863 20806 28868
rect 12998 28573 20511 28863
rect 20801 28573 20806 28863
rect 12998 28568 20806 28573
rect 29480 28218 30980 28238
rect 29480 27918 29560 28218
rect 29550 27858 29560 27918
rect 29960 28148 30980 28218
rect 31283 28148 31461 28153
rect 29960 28147 31462 28148
rect 29960 27969 31283 28147
rect 31461 27969 31462 28147
rect 29960 27968 31462 27969
rect 29960 27918 30980 27968
rect 31283 27963 31461 27968
rect 29960 27858 29970 27918
rect 29550 27853 29970 27858
rect 30530 27143 30750 27148
rect 30530 26933 30535 27143
rect 30745 26933 30750 27143
rect 24740 25238 26600 25318
rect 30530 25278 30750 26933
rect 24740 25078 26380 25238
rect 26540 25078 26600 25238
rect 28360 25218 30750 25278
rect 28360 25098 28400 25218
rect 28540 25098 30750 25218
rect 19991 24208 20289 24213
rect 19990 24207 22150 24208
rect 19990 23909 19991 24207
rect 20289 24203 22150 24207
rect 20289 23913 21855 24203
rect 22145 23913 22150 24203
rect 20289 23909 22150 23913
rect 19990 23908 22150 23909
rect 19991 23903 20289 23908
rect 24760 23538 25000 25078
rect 26370 25073 26550 25078
rect 28360 25058 30750 25098
rect 24760 23298 30500 23538
rect 30740 23298 30746 23538
rect 12998 21025 15296 21030
rect 12998 20735 15001 21025
rect 15291 20735 15296 21025
rect 12998 20730 15296 20735
rect 6431 12990 6729 12995
rect 12998 12990 13298 20730
rect 6430 12989 13298 12990
rect 6430 12691 6431 12989
rect 6729 12691 13298 12989
rect 6430 12690 13298 12691
rect 6431 12685 6729 12690
rect 12998 7070 13298 12690
rect 20895 9210 21193 9215
rect 20894 9209 21878 9210
rect 20894 8911 20895 9209
rect 21193 9205 21878 9209
rect 21193 8915 21583 9205
rect 21873 8915 21878 9205
rect 21193 8911 21878 8915
rect 20894 8910 21878 8911
rect 20895 8905 21193 8910
rect 12998 7065 20806 7070
rect 12998 6775 20511 7065
rect 20801 6775 20806 7065
rect 12998 6770 20806 6775
rect 29480 6420 30980 6440
rect 29480 6120 29560 6420
rect 29550 6060 29560 6120
rect 29960 6350 30980 6420
rect 31283 6350 31461 6355
rect 29960 6349 31462 6350
rect 29960 6171 31283 6349
rect 31461 6171 31462 6349
rect 29960 6170 31462 6171
rect 29960 6120 30980 6170
rect 31283 6165 31461 6170
rect 29960 6060 29970 6120
rect 29550 6055 29970 6060
rect 30530 5345 30750 5350
rect 30530 5135 30535 5345
rect 30745 5135 30750 5345
rect 24740 3440 26600 3520
rect 30530 3480 30750 5135
rect 24740 3280 26380 3440
rect 26540 3280 26600 3440
rect 28360 3420 30750 3480
rect 28360 3300 28400 3420
rect 28540 3300 30750 3420
rect 19991 2410 20289 2415
rect 19990 2409 22150 2410
rect 19990 2111 19991 2409
rect 20289 2405 22150 2409
rect 20289 2115 21855 2405
rect 22145 2115 22150 2405
rect 20289 2111 22150 2115
rect 19990 2110 22150 2111
rect 19991 2105 20289 2110
rect 24760 1740 25000 3280
rect 26370 3275 26550 3280
rect 28360 3260 30750 3300
rect 24760 1500 30500 1740
rect 30740 1500 30746 1740
<< via3 >>
rect 4772 34488 5072 34788
rect 20895 30709 21193 31007
rect 31283 27969 31461 28147
rect 19991 23909 20289 24207
rect 30500 23298 30740 23538
rect 6431 12691 6729 12989
rect 20895 8911 21193 9209
rect 31283 6171 31461 6349
rect 19991 2111 20289 2409
rect 30500 1500 30740 1740
<< metal4 >>
rect 798 44770 858 45152
rect 1534 44770 1594 45152
rect 2270 44770 2330 45152
rect 3006 44770 3066 45152
rect 3742 44770 3802 45152
rect 4478 44770 4538 45152
rect 5214 44770 5274 45152
rect 5950 44770 6010 45152
rect 6686 44770 6746 45152
rect 7422 44770 7482 45152
rect 8158 44770 8218 45152
rect 8894 44770 8954 45152
rect 9630 44770 9690 45152
rect 10366 44770 10426 45152
rect 11102 44770 11162 45152
rect 11838 44770 11898 45152
rect 12574 44770 12634 45152
rect 13310 44770 13370 45152
rect 14046 44770 14106 45152
rect 14782 44770 14842 45152
rect 15518 44770 15578 45152
rect 16254 44770 16314 45152
rect 16990 44770 17050 45152
rect 17726 44770 17786 45152
rect 18462 44952 18522 45152
rect 19198 44952 19258 45152
rect 19934 44952 19994 45152
rect 20670 44952 20730 45152
rect 21406 44952 21466 45152
rect 22142 44952 22202 45152
rect 22878 44952 22938 45152
rect 23614 44952 23674 45152
rect 24350 44952 24410 45152
rect 25086 44952 25146 45152
rect 25822 44952 25882 45152
rect 26558 44952 26618 45152
rect 27294 44952 27354 45152
rect 28030 44952 28090 45152
rect 28766 44952 28826 45152
rect 29502 44952 29562 45152
rect 30238 44952 30298 45152
rect 30974 44952 31034 45152
rect 31710 44952 31770 45152
rect 570 44710 17786 44770
rect 9930 44152 9990 44710
rect 200 34788 500 44152
rect 4771 34788 5073 34789
rect 190 34488 4772 34788
rect 5072 34488 5073 34788
rect 200 12990 500 34488
rect 4771 34487 5073 34488
rect 9800 31008 10100 44152
rect 9800 31007 21194 31008
rect 9800 30709 20895 31007
rect 21193 30709 21194 31007
rect 9800 30708 21194 30709
rect 200 12989 6730 12990
rect 200 12691 6431 12989
rect 6729 12691 6730 12989
rect 200 12690 6730 12691
rect 200 1000 500 12690
rect 9800 9210 10100 30708
rect 19982 28026 20282 30708
rect 31282 28147 31462 28148
rect 19982 27222 20290 28026
rect 19990 24207 20290 27222
rect 19990 23909 19991 24207
rect 20289 23909 20290 24207
rect 19990 23908 20290 23909
rect 31282 27969 31283 28147
rect 31461 27969 31462 28147
rect 30499 23538 30741 23539
rect 31282 23538 31462 27969
rect 30499 23298 30500 23538
rect 30740 23298 31462 23538
rect 30499 23297 30741 23298
rect 9800 9209 21194 9210
rect 9800 8911 20895 9209
rect 21193 8911 21194 9209
rect 9800 8910 21194 8911
rect 9800 1000 10100 8910
rect 19982 6228 20282 8910
rect 31282 8234 31462 23298
rect 23828 8054 31462 8234
rect 19982 5424 20290 6228
rect 19990 2409 20290 5424
rect 19990 2111 19991 2409
rect 20289 2111 20290 2409
rect 19990 2110 20290 2111
rect 23828 926 24008 8054
rect 31282 6349 31462 6350
rect 31282 6171 31283 6349
rect 31461 6171 31462 6349
rect 30499 1740 30741 1741
rect 31282 1740 31462 6171
rect 30499 1500 30500 1740
rect 30740 1500 31462 1740
rect 30499 1499 30741 1500
rect 23828 746 27052 926
rect 370 0 550 200
rect 4786 0 4966 200
rect 9202 0 9382 200
rect 13618 0 13798 200
rect 18034 0 18214 200
rect 22450 0 22630 200
rect 26866 0 27046 746
rect 31282 0 31462 1500
use bandgap  bandgap_0
timestamp 1717066714
transform 1 0 19234 0 1 9074
box -2000 1000 11976 12200
use bandgap_dtmos  bandgap_dtmos_0
timestamp 1717152537
transform 1 0 19234 0 1 30872
box -2000 1000 11977 12200
use p3_opamp  p3_opamp_0
timestamp 1715778954
transform 1 0 21684 0 1 20702
box 3650 3170 8500 8260
use p3_opamp  p3_opamp_1
timestamp 1715778954
transform 1 0 21684 0 1 -1096
box 3650 3170 8500 8260
<< labels >>
flabel metal4 s 30974 44952 31034 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 31710 44952 31770 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 30238 44952 30298 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 31282 0 31462 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26866 0 27046 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22450 0 22630 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18034 0 18214 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 13618 0 13798 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 9202 0 9382 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 4786 0 4966 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 370 0 550 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 29502 44952 29562 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 28030 44952 28090 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 27294 44952 27354 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 25822 44952 25882 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 25086 44952 25146 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23614 44952 23674 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22878 44952 22938 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21406 44952 21466 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 20670 44952 20730 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19198 44952 19258 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 18462 44952 18522 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 5950 44952 6010 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 5214 44952 5274 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 4478 44952 4538 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 3742 44952 3802 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 3006 44952 3066 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 2270 44952 2330 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 1534 44952 1594 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 798 44952 858 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 11838 44952 11898 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 10366 44952 10426 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 9630 44952 9690 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 8158 44952 8218 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 7422 44952 7482 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 16990 44952 17050 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 16254 44952 16314 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 14782 44952 14842 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 14046 44952 14106 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 12574 44952 12634 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 500 44152 1 FreeSans 4800 0 0 0 VPWR
port 51 nsew power bidirectional
flabel metal4 9800 1000 10100 44152 1 FreeSans 4800 0 0 0 VGND
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
