** sch_path: /home/matt/work/asic-workshop/shuttle-2404/tt07-bandgap/xschem/bandgap.sch
.subckt bandgap VDD vref VSS
*.PININFO VSS:B VDD:B vref:B
XM1 top_gate top_gate VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 m=1
XM2 n_gate top_gate VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 m=1
XM3 vref top_gate VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 m=1
XM4 top_gate n_gate Va VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM5 n_gate n_gate Vb VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM6 VSS VSS r4_m6 VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 m=1
XM7 VSS VSS Vb VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 m=1
XM8 VSS VSS r1_m8 VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 m=1
XR4 r4_m6 Va VSS sky130_fd_pr__res_high_po_0p69 L=10 mult=1 m=1
XR1 r1_m8 vref VSS sky130_fd_pr__res_high_po_0p69 L=10 mult=1 m=1
.ends
.end
