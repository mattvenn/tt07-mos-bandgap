magic
tech sky130A
magscale 1 2
timestamp 1712811291
<< nwell >>
rect -1541 -319 1541 319
<< pmoslvt >>
rect -1345 -100 -945 100
rect -887 -100 -487 100
rect -429 -100 -29 100
rect 29 -100 429 100
rect 487 -100 887 100
rect 945 -100 1345 100
<< pdiff >>
rect -1403 88 -1345 100
rect -1403 -88 -1391 88
rect -1357 -88 -1345 88
rect -1403 -100 -1345 -88
rect -945 88 -887 100
rect -945 -88 -933 88
rect -899 -88 -887 88
rect -945 -100 -887 -88
rect -487 88 -429 100
rect -487 -88 -475 88
rect -441 -88 -429 88
rect -487 -100 -429 -88
rect -29 88 29 100
rect -29 -88 -17 88
rect 17 -88 29 88
rect -29 -100 29 -88
rect 429 88 487 100
rect 429 -88 441 88
rect 475 -88 487 88
rect 429 -100 487 -88
rect 887 88 945 100
rect 887 -88 899 88
rect 933 -88 945 88
rect 887 -100 945 -88
rect 1345 88 1403 100
rect 1345 -88 1357 88
rect 1391 -88 1403 88
rect 1345 -100 1403 -88
<< pdiffc >>
rect -1391 -88 -1357 88
rect -933 -88 -899 88
rect -475 -88 -441 88
rect -17 -88 17 88
rect 441 -88 475 88
rect 899 -88 933 88
rect 1357 -88 1391 88
<< nsubdiff >>
rect -1505 249 -1409 283
rect 1409 249 1505 283
rect -1505 187 -1471 249
rect 1471 187 1505 249
rect -1505 -249 -1471 -187
rect 1471 -249 1505 -187
rect -1505 -283 -1409 -249
rect 1409 -283 1505 -249
<< nsubdiffcont >>
rect -1409 249 1409 283
rect -1505 -187 -1471 187
rect 1471 -187 1505 187
rect -1409 -283 1409 -249
<< poly >>
rect -1345 181 -945 197
rect -1345 147 -1329 181
rect -961 147 -945 181
rect -1345 100 -945 147
rect -887 181 -487 197
rect -887 147 -871 181
rect -503 147 -487 181
rect -887 100 -487 147
rect -429 181 -29 197
rect -429 147 -413 181
rect -45 147 -29 181
rect -429 100 -29 147
rect 29 181 429 197
rect 29 147 45 181
rect 413 147 429 181
rect 29 100 429 147
rect 487 181 887 197
rect 487 147 503 181
rect 871 147 887 181
rect 487 100 887 147
rect 945 181 1345 197
rect 945 147 961 181
rect 1329 147 1345 181
rect 945 100 1345 147
rect -1345 -147 -945 -100
rect -1345 -181 -1329 -147
rect -961 -181 -945 -147
rect -1345 -197 -945 -181
rect -887 -147 -487 -100
rect -887 -181 -871 -147
rect -503 -181 -487 -147
rect -887 -197 -487 -181
rect -429 -147 -29 -100
rect -429 -181 -413 -147
rect -45 -181 -29 -147
rect -429 -197 -29 -181
rect 29 -147 429 -100
rect 29 -181 45 -147
rect 413 -181 429 -147
rect 29 -197 429 -181
rect 487 -147 887 -100
rect 487 -181 503 -147
rect 871 -181 887 -147
rect 487 -197 887 -181
rect 945 -147 1345 -100
rect 945 -181 961 -147
rect 1329 -181 1345 -147
rect 945 -197 1345 -181
<< polycont >>
rect -1329 147 -961 181
rect -871 147 -503 181
rect -413 147 -45 181
rect 45 147 413 181
rect 503 147 871 181
rect 961 147 1329 181
rect -1329 -181 -961 -147
rect -871 -181 -503 -147
rect -413 -181 -45 -147
rect 45 -181 413 -147
rect 503 -181 871 -147
rect 961 -181 1329 -147
<< locali >>
rect -1505 249 -1409 283
rect 1409 249 1505 283
rect -1505 187 -1471 249
rect 1471 187 1505 249
rect -1345 147 -1329 181
rect -961 147 -945 181
rect -887 147 -871 181
rect -503 147 -487 181
rect -429 147 -413 181
rect -45 147 -29 181
rect 29 147 45 181
rect 413 147 429 181
rect 487 147 503 181
rect 871 147 887 181
rect 945 147 961 181
rect 1329 147 1345 181
rect -1391 88 -1357 104
rect -1391 -104 -1357 -88
rect -933 88 -899 104
rect -933 -104 -899 -88
rect -475 88 -441 104
rect -475 -104 -441 -88
rect -17 88 17 104
rect -17 -104 17 -88
rect 441 88 475 104
rect 441 -104 475 -88
rect 899 88 933 104
rect 899 -104 933 -88
rect 1357 88 1391 104
rect 1357 -104 1391 -88
rect -1345 -181 -1329 -147
rect -961 -181 -945 -147
rect -887 -181 -871 -147
rect -503 -181 -487 -147
rect -429 -181 -413 -147
rect -45 -181 -29 -147
rect 29 -181 45 -147
rect 413 -181 429 -147
rect 487 -181 503 -147
rect 871 -181 887 -147
rect 945 -181 961 -147
rect 1329 -181 1345 -147
rect -1505 -249 -1471 -187
rect 1471 -249 1505 -187
rect -1505 -283 -1409 -249
rect 1409 -283 1505 -249
<< viali >>
rect -1329 147 -961 181
rect -871 147 -503 181
rect -413 147 -45 181
rect 45 147 413 181
rect 503 147 871 181
rect 961 147 1329 181
rect -1391 -88 -1357 88
rect -933 -88 -899 88
rect -475 -88 -441 88
rect -17 -88 17 88
rect 441 -88 475 88
rect 899 -88 933 88
rect 1357 -88 1391 88
rect -1329 -181 -961 -147
rect -871 -181 -503 -147
rect -413 -181 -45 -147
rect 45 -181 413 -147
rect 503 -181 871 -147
rect 961 -181 1329 -147
<< metal1 >>
rect -1341 181 -949 187
rect -1341 147 -1329 181
rect -961 147 -949 181
rect -1341 141 -949 147
rect -883 181 -491 187
rect -883 147 -871 181
rect -503 147 -491 181
rect -883 141 -491 147
rect -425 181 -33 187
rect -425 147 -413 181
rect -45 147 -33 181
rect -425 141 -33 147
rect 33 181 425 187
rect 33 147 45 181
rect 413 147 425 181
rect 33 141 425 147
rect 491 181 883 187
rect 491 147 503 181
rect 871 147 883 181
rect 491 141 883 147
rect 949 181 1341 187
rect 949 147 961 181
rect 1329 147 1341 181
rect 949 141 1341 147
rect -1397 88 -1351 100
rect -1397 -88 -1391 88
rect -1357 -88 -1351 88
rect -1397 -100 -1351 -88
rect -939 88 -893 100
rect -939 -88 -933 88
rect -899 -88 -893 88
rect -939 -100 -893 -88
rect -481 88 -435 100
rect -481 -88 -475 88
rect -441 -88 -435 88
rect -481 -100 -435 -88
rect -23 88 23 100
rect -23 -88 -17 88
rect 17 -88 23 88
rect -23 -100 23 -88
rect 435 88 481 100
rect 435 -88 441 88
rect 475 -88 481 88
rect 435 -100 481 -88
rect 893 88 939 100
rect 893 -88 899 88
rect 933 -88 939 88
rect 893 -100 939 -88
rect 1351 88 1397 100
rect 1351 -88 1357 88
rect 1391 -88 1397 88
rect 1351 -100 1397 -88
rect -1341 -147 -949 -141
rect -1341 -181 -1329 -147
rect -961 -181 -949 -147
rect -1341 -187 -949 -181
rect -883 -147 -491 -141
rect -883 -181 -871 -147
rect -503 -181 -491 -147
rect -883 -187 -491 -181
rect -425 -147 -33 -141
rect -425 -181 -413 -147
rect -45 -181 -33 -147
rect -425 -187 -33 -181
rect 33 -147 425 -141
rect 33 -181 45 -147
rect 413 -181 425 -147
rect 33 -187 425 -181
rect 491 -147 883 -141
rect 491 -181 503 -147
rect 871 -181 883 -147
rect 491 -187 883 -181
rect 949 -147 1341 -141
rect 949 -181 961 -147
rect 1329 -181 1341 -147
rect 949 -187 1341 -181
<< properties >>
string FIXED_BBOX -1488 -266 1488 266
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 1.0 l 2.0 m 1 nf 6 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
